module tb_task3(output err);
  // your implementation here
endmodule: tb_task3
