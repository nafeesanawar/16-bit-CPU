module tb_task2(output err);
  // your implementation here
endmodule: tb_task2
